package pkg;
        import uvm_pkg::*;
        `include "uvm_macros.svh"
        `include "seq_item.sv"
        `include "sequencer.sv"
        `include "sequence.sv"
        `include "driver.sv"
        `include "monitor.sv"
        `include "agent.sv"
        `include "scoreboard.sv"
		`include "subscriber.sv"
        `include "environment.sv"
        `include "test.sv"
endpackage
